module our;
initial begin $display("hello world"); end
endmodule
